module module2;
endmodule