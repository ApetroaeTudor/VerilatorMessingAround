module pass_through(
    input  wire a,
    output wire y
);
    module2 DUT();
    assign y = a;
endmodule
